module mult_ip (
		input  wire [7:0]  dataa,  //  mult_input.dataa
		input  wire [7:0]  datab,  //            .datab
		input  wire        clock,  //            .clock
		input  wire        aclr,   //            .aclr
		output wire [15:0] result  // mult_output.result
	);
endmodule

